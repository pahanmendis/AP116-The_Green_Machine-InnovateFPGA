// GreenMachine.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module GreenMachine (
		input  wire        clk_clk,                 //               clk.clk
		input  wire        hc05_uart_connect_rxd,   // hc05_uart_connect.rxd
		output wire        hc05_uart_connect_txd,   //                  .txd
		output wire [12:0] memory_mem_a,            //            memory.mem_a
		output wire [2:0]  memory_mem_ba,           //                  .mem_ba
		output wire        memory_mem_ck,           //                  .mem_ck
		output wire        memory_mem_ck_n,         //                  .mem_ck_n
		output wire        memory_mem_cke,          //                  .mem_cke
		output wire        memory_mem_cs_n,         //                  .mem_cs_n
		output wire        memory_mem_ras_n,        //                  .mem_ras_n
		output wire        memory_mem_cas_n,        //                  .mem_cas_n
		output wire        memory_mem_we_n,         //                  .mem_we_n
		output wire        memory_mem_reset_n,      //                  .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,           //                  .mem_dq
		inout  wire        memory_mem_dqs,          //                  .mem_dqs
		inout  wire        memory_mem_dqs_n,        //                  .mem_dqs_n
		output wire        memory_mem_odt,          //                  .mem_odt
		output wire        memory_mem_dm,           //                  .mem_dm
		input  wire        memory_oct_rzqin,        //                  .oct_rzqin
		output wire        mode_control_out_export, //  mode_control_out.export
		input  wire        pio_key_input_export,    //     pio_key_input.export
		input  wire        reset_reset_n            //             reset.reset_n
	);

	wire   [1:0] hps_0_h2f_axi_master_awburst;                     // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                       // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [7:0] hps_0_h2f_axi_master_wstrb;                       // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                      // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                         // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                      // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                       // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                         // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                     // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                      // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                      // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                      // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                      // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [63:0] hps_0_h2f_axi_master_wdata;                       // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                     // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                     // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                        // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                      // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                      // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                      // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                       // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                     // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [63:0] hps_0_h2f_axi_master_rdata;                       // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                     // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                     // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                      // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                      // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                       // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                       // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                       // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                        // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                         // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                      // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                      // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                     // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                      // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect; // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable; // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_hc05_uart_s1_chipselect;        // mm_interconnect_0:hc05_uart_s1_chipselect -> hc05_uart:chipselect
	wire  [15:0] mm_interconnect_0_hc05_uart_s1_readdata;          // hc05_uart:readdata -> mm_interconnect_0:hc05_uart_s1_readdata
	wire   [2:0] mm_interconnect_0_hc05_uart_s1_address;           // mm_interconnect_0:hc05_uart_s1_address -> hc05_uart:address
	wire         mm_interconnect_0_hc05_uart_s1_read;              // mm_interconnect_0:hc05_uart_s1_read -> hc05_uart:read_n
	wire         mm_interconnect_0_hc05_uart_s1_begintransfer;     // mm_interconnect_0:hc05_uart_s1_begintransfer -> hc05_uart:begintransfer
	wire         mm_interconnect_0_hc05_uart_s1_write;             // mm_interconnect_0:hc05_uart_s1_write -> hc05_uart:write_n
	wire  [15:0] mm_interconnect_0_hc05_uart_s1_writedata;         // mm_interconnect_0:hc05_uart_s1_writedata -> hc05_uart:writedata
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                  // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                    // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                    // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                   // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                   // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                    // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                      // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                  // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                   // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                   // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                   // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                   // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                    // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                  // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                  // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                     // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                   // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                   // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                   // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                  // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                   // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                   // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                    // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                     // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                   // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                   // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                  // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                   // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_pio_key_s1_readdata;            // pio_key:readdata -> mm_interconnect_1:pio_key_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_key_s1_address;             // mm_interconnect_1:pio_key_s1_address -> pio_key:address
	wire         mm_interconnect_1_mode_control_s1_chipselect;     // mm_interconnect_1:mode_control_s1_chipselect -> mode_control:chipselect
	wire  [31:0] mm_interconnect_1_mode_control_s1_readdata;       // mode_control:readdata -> mm_interconnect_1:mode_control_s1_readdata
	wire   [1:0] mm_interconnect_1_mode_control_s1_address;        // mm_interconnect_1:mode_control_s1_address -> mode_control:address
	wire         mm_interconnect_1_mode_control_s1_write;          // mm_interconnect_1:mode_control_s1_write -> mode_control:write_n
	wire  [31:0] mm_interconnect_1_mode_control_s1_writedata;      // mm_interconnect_1:mode_control_s1_writedata -> mode_control:writedata
	wire  [31:0] system_console_master_readdata;                   // mm_interconnect_2:system_console_master_readdata -> system_console:master_readdata
	wire         system_console_master_waitrequest;                // mm_interconnect_2:system_console_master_waitrequest -> system_console:master_waitrequest
	wire  [31:0] system_console_master_address;                    // system_console:master_address -> mm_interconnect_2:system_console_master_address
	wire         system_console_master_read;                       // system_console:master_read -> mm_interconnect_2:system_console_master_read
	wire   [3:0] system_console_master_byteenable;                 // system_console:master_byteenable -> mm_interconnect_2:system_console_master_byteenable
	wire         system_console_master_readdatavalid;              // mm_interconnect_2:system_console_master_readdatavalid -> system_console:master_readdatavalid
	wire         system_console_master_write;                      // system_console:master_write -> mm_interconnect_2:system_console_master_write
	wire  [31:0] system_console_master_writedata;                  // system_console:master_writedata -> mm_interconnect_2:system_console_master_writedata
	wire   [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_awburst;    // mm_interconnect_2:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire   [4:0] mm_interconnect_2_hps_0_f2h_axi_slave_awuser;     // mm_interconnect_2:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_arlen;      // mm_interconnect_2:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_wstrb;      // mm_interconnect_2:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_wready;     // hps_0:f2h_WREADY -> mm_interconnect_2:hps_0_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_rid;        // hps_0:f2h_RID -> mm_interconnect_2:hps_0_f2h_axi_slave_rid
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_rready;     // mm_interconnect_2:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire   [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_awlen;      // mm_interconnect_2:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire   [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_wid;        // mm_interconnect_2:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire   [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_arcache;    // mm_interconnect_2:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_wvalid;     // mm_interconnect_2:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire  [31:0] mm_interconnect_2_hps_0_f2h_axi_slave_araddr;     // mm_interconnect_2:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire   [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_arprot;     // mm_interconnect_2:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire   [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_awprot;     // mm_interconnect_2:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [63:0] mm_interconnect_2_hps_0_f2h_axi_slave_wdata;      // mm_interconnect_2:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_arvalid;    // mm_interconnect_2:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire   [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_awcache;    // mm_interconnect_2:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire   [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_arid;       // mm_interconnect_2:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire   [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_arlock;     // mm_interconnect_2:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire   [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_awlock;     // mm_interconnect_2:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire  [31:0] mm_interconnect_2_hps_0_f2h_axi_slave_awaddr;     // mm_interconnect_2:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire   [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_bresp;      // hps_0:f2h_BRESP -> mm_interconnect_2:hps_0_f2h_axi_slave_bresp
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_arready;    // hps_0:f2h_ARREADY -> mm_interconnect_2:hps_0_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_2_hps_0_f2h_axi_slave_rdata;      // hps_0:f2h_RDATA -> mm_interconnect_2:hps_0_f2h_axi_slave_rdata
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_awready;    // hps_0:f2h_AWREADY -> mm_interconnect_2:hps_0_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_arburst;    // mm_interconnect_2:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire   [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_arsize;     // mm_interconnect_2:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_bready;     // mm_interconnect_2:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_rlast;      // hps_0:f2h_RLAST -> mm_interconnect_2:hps_0_f2h_axi_slave_rlast
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_wlast;      // mm_interconnect_2:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire   [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_rresp;      // hps_0:f2h_RRESP -> mm_interconnect_2:hps_0_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_awid;       // mm_interconnect_2:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire   [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_bid;        // hps_0:f2h_BID -> mm_interconnect_2:hps_0_f2h_axi_slave_bid
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_bvalid;     // hps_0:f2h_BVALID -> mm_interconnect_2:hps_0_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_awsize;     // mm_interconnect_2:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_awvalid;    // mm_interconnect_2:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire   [4:0] mm_interconnect_2_hps_0_f2h_axi_slave_aruser;     // mm_interconnect_2:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire         mm_interconnect_2_hps_0_f2h_axi_slave_rvalid;     // hps_0:f2h_RVALID -> mm_interconnect_2:hps_0_f2h_axi_slave_rvalid
	wire         irq_mapper_receiver0_irq;                         // hc05_uart:irq -> irq_mapper:receiver0_irq
	wire  [31:0] hps_0_f2h_irq0_irq;                               // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                               // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [hc05_uart:reset_n, mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:pio_key_reset_reset_bridge_in_reset_reset, mm_interconnect_2:system_console_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:system_console_master_translator_reset_reset_bridge_in_reset_reset, mode_control:reset_n, onchip_memory2_0:reset, pio_key:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;               // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]
	wire         hps_0_h2f_reset_reset;                            // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	GreenMachine_hc05_uart hc05_uart (
		.clk           (clk_clk),                                      //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address       (mm_interconnect_0_hc05_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_hc05_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_hc05_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_hc05_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_hc05_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_hc05_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_hc05_uart_s1_readdata),      //                    .readdata
		.rxd           (hc05_uart_connect_rxd),                        // external_connection.export
		.txd           (hc05_uart_connect_txd),                        //                    .export
		.irq           (irq_mapper_receiver0_irq)                      //                 irq.irq
	);

	GreenMachine_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.h2f_mpu_eventi     (),                                              //    h2f_mpu_events.eventi
		.h2f_mpu_evento     (),                                              //                  .evento
		.h2f_mpu_standbywfe (),                                              //                  .standbywfe
		.h2f_mpu_standbywfi (),                                              //                  .standbywfi
		.mem_a              (memory_mem_a),                                  //            memory.mem_a
		.mem_ba             (memory_mem_ba),                                 //                  .mem_ba
		.mem_ck             (memory_mem_ck),                                 //                  .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                               //                  .mem_ck_n
		.mem_cke            (memory_mem_cke),                                //                  .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                               //                  .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),                              //                  .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                              //                  .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                               //                  .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),                            //                  .mem_reset_n
		.mem_dq             (memory_mem_dq),                                 //                  .mem_dq
		.mem_dqs            (memory_mem_dqs),                                //                  .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                              //                  .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                //                  .mem_odt
		.mem_dm             (memory_mem_dm),                                 //                  .mem_dm
		.oct_rzqin          (memory_oct_rzqin),                              //                  .oct_rzqin
		.h2f_rst_n          (hps_0_h2f_reset_reset),                         //         h2f_reset.reset_n
		.h2f_axi_clk        (clk_clk),                                       //     h2f_axi_clock.clk
		.h2f_AWID           (hps_0_h2f_axi_master_awid),                     //    h2f_axi_master.awid
		.h2f_AWADDR         (hps_0_h2f_axi_master_awaddr),                   //                  .awaddr
		.h2f_AWLEN          (hps_0_h2f_axi_master_awlen),                    //                  .awlen
		.h2f_AWSIZE         (hps_0_h2f_axi_master_awsize),                   //                  .awsize
		.h2f_AWBURST        (hps_0_h2f_axi_master_awburst),                  //                  .awburst
		.h2f_AWLOCK         (hps_0_h2f_axi_master_awlock),                   //                  .awlock
		.h2f_AWCACHE        (hps_0_h2f_axi_master_awcache),                  //                  .awcache
		.h2f_AWPROT         (hps_0_h2f_axi_master_awprot),                   //                  .awprot
		.h2f_AWVALID        (hps_0_h2f_axi_master_awvalid),                  //                  .awvalid
		.h2f_AWREADY        (hps_0_h2f_axi_master_awready),                  //                  .awready
		.h2f_WID            (hps_0_h2f_axi_master_wid),                      //                  .wid
		.h2f_WDATA          (hps_0_h2f_axi_master_wdata),                    //                  .wdata
		.h2f_WSTRB          (hps_0_h2f_axi_master_wstrb),                    //                  .wstrb
		.h2f_WLAST          (hps_0_h2f_axi_master_wlast),                    //                  .wlast
		.h2f_WVALID         (hps_0_h2f_axi_master_wvalid),                   //                  .wvalid
		.h2f_WREADY         (hps_0_h2f_axi_master_wready),                   //                  .wready
		.h2f_BID            (hps_0_h2f_axi_master_bid),                      //                  .bid
		.h2f_BRESP          (hps_0_h2f_axi_master_bresp),                    //                  .bresp
		.h2f_BVALID         (hps_0_h2f_axi_master_bvalid),                   //                  .bvalid
		.h2f_BREADY         (hps_0_h2f_axi_master_bready),                   //                  .bready
		.h2f_ARID           (hps_0_h2f_axi_master_arid),                     //                  .arid
		.h2f_ARADDR         (hps_0_h2f_axi_master_araddr),                   //                  .araddr
		.h2f_ARLEN          (hps_0_h2f_axi_master_arlen),                    //                  .arlen
		.h2f_ARSIZE         (hps_0_h2f_axi_master_arsize),                   //                  .arsize
		.h2f_ARBURST        (hps_0_h2f_axi_master_arburst),                  //                  .arburst
		.h2f_ARLOCK         (hps_0_h2f_axi_master_arlock),                   //                  .arlock
		.h2f_ARCACHE        (hps_0_h2f_axi_master_arcache),                  //                  .arcache
		.h2f_ARPROT         (hps_0_h2f_axi_master_arprot),                   //                  .arprot
		.h2f_ARVALID        (hps_0_h2f_axi_master_arvalid),                  //                  .arvalid
		.h2f_ARREADY        (hps_0_h2f_axi_master_arready),                  //                  .arready
		.h2f_RID            (hps_0_h2f_axi_master_rid),                      //                  .rid
		.h2f_RDATA          (hps_0_h2f_axi_master_rdata),                    //                  .rdata
		.h2f_RRESP          (hps_0_h2f_axi_master_rresp),                    //                  .rresp
		.h2f_RLAST          (hps_0_h2f_axi_master_rlast),                    //                  .rlast
		.h2f_RVALID         (hps_0_h2f_axi_master_rvalid),                   //                  .rvalid
		.h2f_RREADY         (hps_0_h2f_axi_master_rready),                   //                  .rready
		.f2h_axi_clk        (clk_clk),                                       //     f2h_axi_clock.clk
		.f2h_AWID           (mm_interconnect_2_hps_0_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR         (mm_interconnect_2_hps_0_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN          (mm_interconnect_2_hps_0_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE         (mm_interconnect_2_hps_0_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST        (mm_interconnect_2_hps_0_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK         (mm_interconnect_2_hps_0_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE        (mm_interconnect_2_hps_0_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT         (mm_interconnect_2_hps_0_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID        (mm_interconnect_2_hps_0_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY        (mm_interconnect_2_hps_0_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER         (mm_interconnect_2_hps_0_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID            (mm_interconnect_2_hps_0_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA          (mm_interconnect_2_hps_0_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB          (mm_interconnect_2_hps_0_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST          (mm_interconnect_2_hps_0_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID         (mm_interconnect_2_hps_0_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY         (mm_interconnect_2_hps_0_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID            (mm_interconnect_2_hps_0_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP          (mm_interconnect_2_hps_0_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID         (mm_interconnect_2_hps_0_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY         (mm_interconnect_2_hps_0_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID           (mm_interconnect_2_hps_0_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR         (mm_interconnect_2_hps_0_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN          (mm_interconnect_2_hps_0_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE         (mm_interconnect_2_hps_0_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST        (mm_interconnect_2_hps_0_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK         (mm_interconnect_2_hps_0_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE        (mm_interconnect_2_hps_0_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT         (mm_interconnect_2_hps_0_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID        (mm_interconnect_2_hps_0_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY        (mm_interconnect_2_hps_0_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER         (mm_interconnect_2_hps_0_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID            (mm_interconnect_2_hps_0_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA          (mm_interconnect_2_hps_0_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP          (mm_interconnect_2_hps_0_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST          (mm_interconnect_2_hps_0_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID         (mm_interconnect_2_hps_0_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY         (mm_interconnect_2_hps_0_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk     (clk_clk),                                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID        (hps_0_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR      (hps_0_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN       (hps_0_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE      (hps_0_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST     (hps_0_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK      (hps_0_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE     (hps_0_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT      (hps_0_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID     (hps_0_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY     (hps_0_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID         (hps_0_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA       (hps_0_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB       (hps_0_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST       (hps_0_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID      (hps_0_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY      (hps_0_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID         (hps_0_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP       (hps_0_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID      (hps_0_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY      (hps_0_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID        (hps_0_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR      (hps_0_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN       (hps_0_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE      (hps_0_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST     (hps_0_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK      (hps_0_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE     (hps_0_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT      (hps_0_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID     (hps_0_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY     (hps_0_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID         (hps_0_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA       (hps_0_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP       (hps_0_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST       (hps_0_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID      (hps_0_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY      (hps_0_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0         (hps_0_f2h_irq0_irq),                            //          f2h_irq0.irq
		.f2h_irq_p1         (hps_0_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	GreenMachine_mode_control mode_control (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_mode_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_mode_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_mode_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_mode_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_mode_control_s1_readdata),   //                    .readdata
		.out_port   (mode_control_out_export)                       // external_connection.export
	);

	GreenMachine_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	GreenMachine_pio_key pio_key (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_1_pio_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_pio_key_s1_readdata), //                    .readdata
		.in_port  (pio_key_input_export)                   // external_connection.export
	);

	GreenMachine_system_console #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) system_console (
		.clk_clk              (clk_clk),                             //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                      //    clk_reset.reset
		.master_address       (system_console_master_address),       //       master.address
		.master_readdata      (system_console_master_readdata),      //             .readdata
		.master_read          (system_console_master_read),          //             .read
		.master_write         (system_console_master_write),         //             .write
		.master_writedata     (system_console_master_writedata),     //             .writedata
		.master_waitrequest   (system_console_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (system_console_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (system_console_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                     // master_reset.reset
	);

	GreenMachine_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                        //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                      //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                       //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                      //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                     //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                      //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                     //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                      //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                     //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                     //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                         //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                       //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                       //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                       //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                      //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                      //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                         //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                       //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                      //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                      //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                        //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                      //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                       //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                      //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                     //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                      //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                     //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                      //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                     //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                     //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                         //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                       //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                       //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                       //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                      //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                      //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                          //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),               // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                   //              onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.hc05_uart_s1_address                                             (mm_interconnect_0_hc05_uart_s1_address),           //                                               hc05_uart_s1.address
		.hc05_uart_s1_write                                               (mm_interconnect_0_hc05_uart_s1_write),             //                                                           .write
		.hc05_uart_s1_read                                                (mm_interconnect_0_hc05_uart_s1_read),              //                                                           .read
		.hc05_uart_s1_readdata                                            (mm_interconnect_0_hc05_uart_s1_readdata),          //                                                           .readdata
		.hc05_uart_s1_writedata                                           (mm_interconnect_0_hc05_uart_s1_writedata),         //                                                           .writedata
		.hc05_uart_s1_begintransfer                                       (mm_interconnect_0_hc05_uart_s1_begintransfer),     //                                                           .begintransfer
		.hc05_uart_s1_chipselect                                          (mm_interconnect_0_hc05_uart_s1_chipselect),        //                                                           .chipselect
		.onchip_memory2_0_s1_address                                      (mm_interconnect_0_onchip_memory2_0_s1_address),    //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                                           .clken
	);

	GreenMachine_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                 //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),               //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),               //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),              //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),               //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),              //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),               //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),              //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),              //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                  //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),               //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),               //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                  //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),               //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),               //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                 //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),               //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),               //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),              //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),               //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),              //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),               //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),              //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),              //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                  //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),               //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),               //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                      //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),           // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pio_key_reset_reset_bridge_in_reset_reset                           (rst_controller_reset_out_reset),               //                           pio_key_reset_reset_bridge_in_reset.reset
		.mode_control_s1_address                                             (mm_interconnect_1_mode_control_s1_address),    //                                               mode_control_s1.address
		.mode_control_s1_write                                               (mm_interconnect_1_mode_control_s1_write),      //                                                              .write
		.mode_control_s1_readdata                                            (mm_interconnect_1_mode_control_s1_readdata),   //                                                              .readdata
		.mode_control_s1_writedata                                           (mm_interconnect_1_mode_control_s1_writedata),  //                                                              .writedata
		.mode_control_s1_chipselect                                          (mm_interconnect_1_mode_control_s1_chipselect), //                                                              .chipselect
		.pio_key_s1_address                                                  (mm_interconnect_1_pio_key_s1_address),         //                                                    pio_key_s1.address
		.pio_key_s1_readdata                                                 (mm_interconnect_1_pio_key_s1_readdata)         //                                                              .readdata
	);

	GreenMachine_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_f2h_axi_slave_awid                                           (mm_interconnect_2_hps_0_f2h_axi_slave_awid),    //                                          hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awaddr),  //                                                             .awaddr
		.hps_0_f2h_axi_slave_awlen                                          (mm_interconnect_2_hps_0_f2h_axi_slave_awlen),   //                                                             .awlen
		.hps_0_f2h_axi_slave_awsize                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awsize),  //                                                             .awsize
		.hps_0_f2h_axi_slave_awburst                                        (mm_interconnect_2_hps_0_f2h_axi_slave_awburst), //                                                             .awburst
		.hps_0_f2h_axi_slave_awlock                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awlock),  //                                                             .awlock
		.hps_0_f2h_axi_slave_awcache                                        (mm_interconnect_2_hps_0_f2h_axi_slave_awcache), //                                                             .awcache
		.hps_0_f2h_axi_slave_awprot                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awprot),  //                                                             .awprot
		.hps_0_f2h_axi_slave_awuser                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awuser),  //                                                             .awuser
		.hps_0_f2h_axi_slave_awvalid                                        (mm_interconnect_2_hps_0_f2h_axi_slave_awvalid), //                                                             .awvalid
		.hps_0_f2h_axi_slave_awready                                        (mm_interconnect_2_hps_0_f2h_axi_slave_awready), //                                                             .awready
		.hps_0_f2h_axi_slave_wid                                            (mm_interconnect_2_hps_0_f2h_axi_slave_wid),     //                                                             .wid
		.hps_0_f2h_axi_slave_wdata                                          (mm_interconnect_2_hps_0_f2h_axi_slave_wdata),   //                                                             .wdata
		.hps_0_f2h_axi_slave_wstrb                                          (mm_interconnect_2_hps_0_f2h_axi_slave_wstrb),   //                                                             .wstrb
		.hps_0_f2h_axi_slave_wlast                                          (mm_interconnect_2_hps_0_f2h_axi_slave_wlast),   //                                                             .wlast
		.hps_0_f2h_axi_slave_wvalid                                         (mm_interconnect_2_hps_0_f2h_axi_slave_wvalid),  //                                                             .wvalid
		.hps_0_f2h_axi_slave_wready                                         (mm_interconnect_2_hps_0_f2h_axi_slave_wready),  //                                                             .wready
		.hps_0_f2h_axi_slave_bid                                            (mm_interconnect_2_hps_0_f2h_axi_slave_bid),     //                                                             .bid
		.hps_0_f2h_axi_slave_bresp                                          (mm_interconnect_2_hps_0_f2h_axi_slave_bresp),   //                                                             .bresp
		.hps_0_f2h_axi_slave_bvalid                                         (mm_interconnect_2_hps_0_f2h_axi_slave_bvalid),  //                                                             .bvalid
		.hps_0_f2h_axi_slave_bready                                         (mm_interconnect_2_hps_0_f2h_axi_slave_bready),  //                                                             .bready
		.hps_0_f2h_axi_slave_arid                                           (mm_interconnect_2_hps_0_f2h_axi_slave_arid),    //                                                             .arid
		.hps_0_f2h_axi_slave_araddr                                         (mm_interconnect_2_hps_0_f2h_axi_slave_araddr),  //                                                             .araddr
		.hps_0_f2h_axi_slave_arlen                                          (mm_interconnect_2_hps_0_f2h_axi_slave_arlen),   //                                                             .arlen
		.hps_0_f2h_axi_slave_arsize                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arsize),  //                                                             .arsize
		.hps_0_f2h_axi_slave_arburst                                        (mm_interconnect_2_hps_0_f2h_axi_slave_arburst), //                                                             .arburst
		.hps_0_f2h_axi_slave_arlock                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arlock),  //                                                             .arlock
		.hps_0_f2h_axi_slave_arcache                                        (mm_interconnect_2_hps_0_f2h_axi_slave_arcache), //                                                             .arcache
		.hps_0_f2h_axi_slave_arprot                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arprot),  //                                                             .arprot
		.hps_0_f2h_axi_slave_aruser                                         (mm_interconnect_2_hps_0_f2h_axi_slave_aruser),  //                                                             .aruser
		.hps_0_f2h_axi_slave_arvalid                                        (mm_interconnect_2_hps_0_f2h_axi_slave_arvalid), //                                                             .arvalid
		.hps_0_f2h_axi_slave_arready                                        (mm_interconnect_2_hps_0_f2h_axi_slave_arready), //                                                             .arready
		.hps_0_f2h_axi_slave_rid                                            (mm_interconnect_2_hps_0_f2h_axi_slave_rid),     //                                                             .rid
		.hps_0_f2h_axi_slave_rdata                                          (mm_interconnect_2_hps_0_f2h_axi_slave_rdata),   //                                                             .rdata
		.hps_0_f2h_axi_slave_rresp                                          (mm_interconnect_2_hps_0_f2h_axi_slave_rresp),   //                                                             .rresp
		.hps_0_f2h_axi_slave_rlast                                          (mm_interconnect_2_hps_0_f2h_axi_slave_rlast),   //                                                             .rlast
		.hps_0_f2h_axi_slave_rvalid                                         (mm_interconnect_2_hps_0_f2h_axi_slave_rvalid),  //                                                             .rvalid
		.hps_0_f2h_axi_slave_rready                                         (mm_interconnect_2_hps_0_f2h_axi_slave_rready),  //                                                             .rready
		.clk_0_clk_clk                                                      (clk_clk),                                       //                                                    clk_0_clk.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),            //   hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.system_console_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                //               system_console_clk_reset_reset_bridge_in_reset.reset
		.system_console_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // system_console_master_translator_reset_reset_bridge_in_reset.reset
		.system_console_master_address                                      (system_console_master_address),                 //                                        system_console_master.address
		.system_console_master_waitrequest                                  (system_console_master_waitrequest),             //                                                             .waitrequest
		.system_console_master_byteenable                                   (system_console_master_byteenable),              //                                                             .byteenable
		.system_console_master_read                                         (system_console_master_read),                    //                                                             .read
		.system_console_master_readdata                                     (system_console_master_readdata),                //                                                             .readdata
		.system_console_master_readdatavalid                                (system_console_master_readdatavalid),           //                                                             .readdatavalid
		.system_console_master_write                                        (system_console_master_write),                   //                                                             .write
		.system_console_master_writedata                                    (system_console_master_writedata)                //                                                             .writedata
	);

	GreenMachine_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	GreenMachine_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
